module AND_gate(IN1,IN2,OUT1);
input IN1,IN2;
output OUT1;

assign OUT1 = IN1 & IN2;

endmodule
